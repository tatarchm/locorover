PK   {n<VB�D  z�     cirkitFile.json�]�s7��W��]9,<�n�fS��n\�Wك�bg01keR�G�����CJ�<@6�[r��-�F�C?��ɦ�ͯ��z����v�^MN>��sq�)�N���n=�uS<~��}�g�?}V�?=�W~���R�[�Y��L9%��]&KV�.�|!�lr���ttw��.p�%��
�O�_T�uX�yel�r]d�5>S��3��EVp�J�L�z��z�\#W��s��\w���B�y�=G��+d��G��#�Ǒ�H�	��E�O �'�j��[��6���\�?S��uQ�5+��T�*3���QC穡Mm��r����y�9_!xiy�͵�{3�A���4¢Ɩ��jl�$r���.�S�`,�+΂�`�l!T����
�Ю���O=1s��32K�̄~�}&��ʔ�eX=k3Uˢ���9�vhdԜ����.��5ό�2S����%��r�(U�e^..���i���@A��Zq��@��6���i�	�vހ(^6��B������9�/����EP����yz���#wx�`,0fl�ۢ�Ny�P�3vj�B=M�������D��r�h�g�n�ˁ���2`9����],6G�$=�2$`k�O�kk�dSW��3�Ի9�ۧ��#́�,��2`9���p�X���.��;2#T2�] 0x��K��oz��R�C/=B
���%�GH�יh�_ʮ���ĀV�ߋ�R�@7]	��\.��� <�?���к0A�E�pQ�Kne%.:r�k�
�����Ȑp�$\��K�^N_N�_�h�h64�4�4 �4(4(D:�łŢA��u��M�b���[���Ιp�M�����6G�ڕ6�KaKWc�.��UCˡ�y��8���6�,^��-SF�x�����Z�a.����ՅV/s�/�.�0x�IC�|3���%?.��U�˨�V�ft�hC�s\�{��jqM���o�
��vټ��b��-��5�ģ�\�8#��ã�_4%��R�D	�<�0F#��	��W�H��s��H4mZNň�lب�D	{8��D#Q¶�*?iH2�Mŉ%�����Ld���K&�ƕ��d"ҹ��K��ƕ��d"S��3��:��t>�`u9��=]�iA�H�nĩ��;����~�)�� <A�E�pQ$\4	����!�bI�8�������������ÜĜłłHӠXРXРXРXРXРXРXРXҠX^E1���rUp=��,�z��UY�� <Y�*=p=���׃�\�*<p=�媺׃PG^�^�<�� 64 ��y��Al�Ճq*F,���ՃH$J q\=�D���ՃH$Jl�q� �;m\=�D"�M˩��W"�(a�ՃH$J��q� I���8���Y���LqSqbIwdd=�F&2�Mŉ%��� �����!���r�]�փ�\�1�u~�}w�4_V�O��N>/7~;|(J_͗��zS������M(`䏩?|�b�Y��aFƜK橑��#L��sB7O��#�a��s�y��u&��5���阱SoA�e�0�sC���9�p�AU
Pcc�y��%��zj��;N�o�!Bڸ��D�v�d�]u����v��%:��B)fh�v	��ÓϺ�ֿ��XUC��� �7sb?����JoH��k8�x�>�E^õ����/
�:�6^��M ��&�}�E@:�x}����*8�9ѫ*�5b�
���Nk��G"*J�$"��C�`�D��"�ؠ�@l숄#�b?`�jD�e���2�zHM"2���)_#��K���c��|�\=_!z�{]_*���v�s��_ �Kd�X�e���t�]"��+��� �[d�E�X|r,@9��9�e��!��c�ȱHX$
���"Q`�(�ʒ#Mm���ty_�&R7�k@~9.���C���I,����ou&�KD��a��a�}�\�]"��J�=��P�?��l��׆`P ��������p,����a|3��|g����	�'�b ��~U��/� ���K�B��?T��磎�?�b��,X_��-����/��BJ�Ӻ�n!����	ճ�u��8�za�[A��E��{�h� �=�6��R��ew���T+�0�#��`� P�xl 95��V�B�<�@�l����R�|#璅��(M����tإ�M�e����:���,�Xn	����ɇį�S�r�`-FXѧ�~x����W4:�Z43hJ�Mq�)o7f�y���=D�!ޱ��=D�!b{4��T�A��@�l���>9�:@2���C���']�8& �1�=�pX�]D���_ !�u�'�[�Q�A{¤���U.]��/�F��	����W�<�O`�A�'�g0⠯��qзN���Ձ�::��Io.��|�">��Jw.<i^�H�KBH�=�r���x��X��h@;O?����DU�i��&�o�&�o��&�oR�&�o��&�oʏMy���L���l���\��?��/^����a~�W��z=Xnw�ת.M]�����LIUeNq�-l��1�r�˹���f��r���]p�����a��p�̝�X�[����7�_?�"@S�������P�0�棷����얾q�?=���a����r�kX�U�)�[��ߊ�}��矾ϸ�Mef�Z�IL�oۏ��?��8O��(hh���/��r���?���_M�va����T��uQ����$�9�I�w���_?�W�ėY����r��4|f������d3���	�6�n�M`1Q����2�ږ/�˪ZTY���"�Q�EЇ�jW��CP|2��7�����d�#\��|��G�^:1�S��00��33�;&��D�d��T:�����ܽ��������3>ca��2 ���݌k��q��R#
PA��eD��A���jcD�ϟ@�
��	�50���z�_���fU�c�0j�d�}�WY�����i���*l�stOċ���` dV�Ȍ�:<nÍ.�Q�����c���F��-�b�M�PC�f�)��Q��x���7��)t�?��^�w�0Q2t�k����S�8{T"��_�1�6 6wA)�u��H)}��!�T%w��ƸL��>TA�>���,�|E=���
n�a�ۢ�L� x~�{���3a�RG��D$����
��N��3-]�u'2�Dg��c�|�LZ1s�*�|�fB0)��]�y'7�A8޴���xа�%�/l+�vg39<I ����L�"Y��|���+rN B����<����Z7�jm�0�����d�	��z��Y��O��;\e W�`u����yh���4��Z1��Yf+���Ef2||�DWK�R� [`�5ػf�\~I�A�z�N�Ԡ��s�=7�߭� x�A$�*�C���C���ms�O��6��
,Z������ �dZ��r7��`�8���Q3'��L6i�}:�t}@ӹ�p4Lׇ�0]e�t膛z&�Ar���5����#�:D$�b�"g"�J�s�dʧ�fȕ|��R�kq^Ȃ��g>h����e�E��R��8YH�}�׃��`Z\O-{��B�������?u�OKv���U�E&Cl|Q1}�ޯ�I�uX�Iƙ����l"��r6CN�|����"���	���o�ػ�3r&%ˣ��{��m��@^�}��s
����v�����_�x_�'�{/�'w�O_~?��������M�4���4�����
V9mXm���(E��F'��z�ڽ-v^_���'1c�S�66�k6�6~z�>��$����\�3�ۧD�<�==G.p"�:�}�z?�����[�)A��@��A�HA�ǀ����?'>����?��r:D@PԵ�L A;: �$7� ����&�yzJ!�R*�A
D%�����[8l�-�T�����t-%�`�vB�d`st�t����Q����[ �P9=X�c.�MuX��]�sPQB�N��b;����t5��$@��"������w�����۩ēb1)k�P`�A���!R�#�K:�֮$��$����������P+ٜ�jи���9�@TP��P�Q�"����������P���jX���QA!T�L��B�B7�^�G�Q�WB�RU@�a���ZD�Pne%!4�,��l����t�v����`)�`�v��7�)����A�%s����D���D���7D��K"��*ĉa�ȶB��a��7S�K�2�F�Q0_
v�����u��(�NB�t)��0���C��L������8Տ4��T`��BvQ�%�I��F%d{�Lh�.���l��@2�ɚ#$�RAu��m�-44 ]�!�nH�� Y`0
j��5r��}��h�MGc]�ID�D��Tи�ٺ����b!���p�d#��(��t�d��B��f�(�(&��	�d��T)�ųˇ���;�Y��]޶�c�_��X틇�ן����m\�_'_�PK   {n<VB�D  z�             ��    cirkitFile.jsonPK      =   4    