PK   :n<V>Y0[�  (�     cirkitFile.json��s�6���{5�@ ����L�d�����h(�9U$/E%�f��hK����Ф��������}B>Fu��nW�������W�mt��"z���Cv�i����٭~��Ǉ���;n�x�q�{����m�9��ik��X��5+M��He��VIts{�����h�9��pݧ:sU�"O���6:�ccs�kVX�S���	#K�Ȝ2rJ[2E�i�V*�D�wF�	bI�O���cD��? �TkK����? �)��:�)c+�؂4�&�M�7`Hc��,'>o|�y�Y"
H��,X�T��Dg"��Z�XK��V��3W��QFNfFN@�][�,+b6w��u,J��|mL",��0�ȤkNgFVzPJ+cy,l^���$���:��i��C���S��]�׍�0�܊#��0322�'��)#��y�y"���#�j��s^�TF��Q���ET��h�t͛\�]a����}�ؤ���;�����8�2��S��o)c��٧��R���jbi)�6i"R�)����"�Z2�,A��Z�LC���A�HѢ�h1a�ozY|Y~��F�Qa�ab�bC1��a(�0C�!��R\�	�������%(�:�ui(�Z�sй))^7��*�آN���nqfV[�qs�"�شl��Cce-ݺȒ�i-�"�����B.k��D.�.��q�NcK��=l��r��-!X]y�:lU�2u�?�]u��|?���':����pt>١�S����e_v���y�Oy��K͛����ن�7ӵ@-<�D��%�EѢ�h1a�ozY|Y~Y�Y�Y�Y�Y�Y�!�����Pa(�0C�!��bC1C1�J1:o�k�:t�L�ru.輙���\�y3]K��\5z輙���C��t-W:o�k�j��ys �����'>o�&��#O|������[�{s|ۼ��ߣ�.�Um���M��b���]]�:���|9����<�~A��G񚔑)un672��R�$edJ�7�o�el�Q����6$�D[��elA�((�5'տ��5��}@Hilʂ���H[�Iy-ilIK���<ym���;W�m�)�~�f��\������������
|��>b�qq_"�O�w\���	?�S G!�@FL��Ч@M����̛d�%P�2^5�_"R"� )Z��i�V�d�L�;� S �P*T|@�L�C�5�0rD�c�.��y���߻�ۤ������eE�B�����ߗL���Lh��v2P7,���P�N�kbC���'�OF�Q	m��$����!�rȨ 2*�@%Ȗ�J"PI*�@%��2��3i~C�@_J�2�G
�X%��T�����CD+*��Q�i1PG���@�Lx��C2����#3���Fp���@�C��d��R$��H������%�k82��L(Ww�����P�_�3��IH
&�Ԗ��3���d�o�S�7���
����":u�
� ;�{�!c��?��� o����	�����3�F�[�
zɶ��>��C��3/μ<������}�=�� �|������"{[����(wx����P��뀹1AW�[q8�խm�M]?�҉\�}<cI:����g�3H��v��=�� ���s'��J۩1\H_�6o���h?�~����rH��1v����>�>�v�%�l}�ύ����v���`�>���m��e�º&6n��	�M�k��&�5�q����ItMb�$�&9nJ��tܤ�&�C�l�Y�k��]V�-2�n�����w�(sU�¹�|.���Z�*��*㫔�`���`���jc�ƣ0���,&���5���c�ћz�h릲m���q���｛쾩���B��;��o]D��������c�y����&r��v^o��4G7e��[׸��/վZo��g��m�4��z�˶�2˛Cm�KS8;���cV���a`*�뽻}մǯ�rŖJ*F�\�<Yj�$ȎV�����r*"�s�l�c-u�ܚ�(��)縸����ɶ��*�[D��r�/;�,j︻�U�olwKo���\p�4�?�~q+���I �.�I�D*��QJ��MN�oU�9�C�#�dK����#�@&eCd3K&�P�J��&�
�QĤ�#���m*��p��$_�����k��]����j�y�-����Ќ�Γ.��{��t��t)�p��9�X[X�"�D�8�Y+ť�݊)�Y%T>����8<�؈�$e��.��L5����g�������~~�$[�Ï?�ֻ&8&������r�X&B+�;#����<K���r���8�����M[�9��Ȇ�R�!%u���؈��e����p��pv�t3�K7m��s��2*���� ��t�}�.A!:���p�ˤB�~���Rr㞺��pz| Ȓ�o:)�5,��J��w1� �\��!M�tR����E�;ǜ�u-��܃��Isv%'�����n4H�f Ƌ9�񬇃<_�s�* �]�X�8��yu�P =j��{�E_��m�Z=L�.��b�����w�R����q�Np����Gj!ڛv��Hx��"᱒2��H�8K`�5w���EZ	T��K&��:�>王�ϝ#�i��|�C<5H�t���������`fs=�i<P���u_�~���ť7`����3=���%��i�6���N�y�I��&��wgZnĴ�a0)7�Ѵ��i�1e�r-t�M#��FHN�]���;l��r7;g袘%z�X*}���G�g��r)��6>TE��U$�,]%|}���Q�Md_��1��������_e��-�.���m���Ke?��UɗZ>�E�����# �ŝ3�Yݼ�������i�2�-.�½XhU�ه�!����3��wնy�5���www��@�.��������Oon��r�3R+.���	!y�z����L��N����>9��PO�	E
�$(�s��W�V�e*y~+B����F�@	��PL$�7k((p/��P�`j(^0�Bі�Nw�%KS�b %ʠ��87KH���a?��J�����=35$d8w�{�2�;z��^
Y���:+~� H��Z��W_�X���C�s4Q /��A�_��J!�=[�Ur����]%���ٽ4~:���m:����'I�ґ�O,Zj�*�z�"Ŵ�D���_*�c\�֞�F�#�Q���Tν�NJL�s�#)��$��~�b),��s��f�i:��c7��٫B��%�3Լ9����R��A/�@J�++��?S=(B�+���������^�����/��w�J
���<����������^�����/��'�E��o)EHD�Y�K&���K��^�����/��	'5��Pm6�˟���U��G7��}�G�?[��m���ݻW�}��k�u��ӟPK   :n<V>Y0[�  (�             ��    cirkitFile.jsonPK      =   �    